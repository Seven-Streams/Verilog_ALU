`include "Add.v"

module Mul(
        input [31:0] a,
        input [31:0] b,
        output [63:0] product
    );
endmodule
